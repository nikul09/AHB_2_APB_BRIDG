`ifndef defines
`define defines

//`define ADDR_WIDTH 32
//`define DATA_WIDTH 32

//typedef enum bit{RD_REQ,WR_REQ}wr_rd_kind;
//typedef enum bit[1:0]{OKAY,ERROR,RETRY,SPLIT}resp_kind;
//typedef enum bit[2:0]{SINGLE,INCR,WRAP4,INCR4,WRAP8,INCR8,WRAP16,INCR16}hbrust_kind;
//typedef enum bit[1:0]{IDLE,BUSY,NONSEQ,SEQ}htrans_kind;

//`define MDRV_CB vinf.m_drv
//`define SMON_CB vinf.s_mon
//`define MMON_CB vinf.m_mon

`endif
